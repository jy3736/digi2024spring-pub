module dff_ne_ar(
    input wire clk,
    input wire rst,
    input wire d,
    output reg q
);

// add your code here

endmodule
