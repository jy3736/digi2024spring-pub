module comb_logic(
    input wire a,
    input wire b,
    input wire c,
    input wire d,
    output reg x,
    output reg y
);

// ======================
// = add your code here =
// ======================

endmodule
