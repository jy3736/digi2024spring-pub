module mux2(input in0, input in1, input sel, output out);
    assign out = sel ? in1 : in0;
endmodule

module hadd(
    input a, b,
    output sum, co);

// ======================
// = add your code here =
// ======================

endmodule

