module hadd(
    input a,
    input b,
    output s,
    output c
);

assign s = a ^ b;
assign c = a & b;

endmodule

module fadd(
    input a,
    input b,
    input cin,
    output s,
    output cout
);

// ======================
// = add your code here =
// ======================

endmodule
