module comb_logic(
    input a,
    input b,
    input c,
    input d,
    output reg x,
    output reg y
);

// add your code here

endmodule
