module shift_register(
    input wire clk,
    input wire rst,
    input wire L,        // Parallel load input
    input wire r0,       // Load/shift control for Q0
    input wire r1,       // Load/shift control for Q1
    input wire r2,       // Load/shift control for Q2
    output reg Q0,
    output reg Q1,
    output reg Q2
);

// add your code here

endmodule
