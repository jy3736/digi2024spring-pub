module dual_edge_dff_ar(
    input wire clk,
    input wire rst,
    input wire d0,
    input wire d1,
    output reg q
);

// add your code here

endmodule
