module filter_logic(
    input a,
    input b,
    input c,
    input d,
    input e,
    input f,
    output reg x,
    output reg y,
    output reg z
);

// add your code here

endmodule
