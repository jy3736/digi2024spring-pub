module mux2(input in0, input in1, input sel, output out);
    assign out = sel ? in1 : in0;
endmodule

module and3(
    input a, b, c,
    output y);
    wire ab;

// ======================
// = add your code here =
// ======================

endmodule
