module comb01(
    input a,
    input b,
    output reg not_a,
    output reg not_b,
    output reg and_ab,
    output reg or_ab,
    output reg xor_ab,
    output reg nand_ab,
    output reg nor_ab,
    output reg xnor_ab
);

// add your code here

endmodule
